module INV(output[15:0] y,input[15:0] x);
  
 
  
 assign y= ~x;
  
  
endmodule  